-- --------------------------------------------------------
-- Hardware software codesign
-- --------------------------------------------------------
-- Course assignments
--
-- File: hamming_distance.vhd (vhdl)
-- By: Lowie Deferme (UHasselt/KULeuven - FIIW)
-- On: 26 February 2022

